module adder (input [31:0] data1, [31:0] data2, output [31:0] out_data);
    assign out_data = data1 + data2;
    
endmodule
